package hs_npu_pkg;
endpackage : hs_npu_pkg
