package hs_npu_pkg;

  typedef logic signed [31:0] word;
  typedef logic signed [15:0] short;
  typedef logic [31:0] uword;


endpackage : hs_npu_pkg
